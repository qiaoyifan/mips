/*
* 将32位数据译码为64位字型码
*/

module Seg8BCD(
		input [31:0] in,
		output reg [63:0] out);


	
	

	always @( * ) begin
		
			
			case(in[3:0])
				4'b0000:out[7:0]=8'b00000011;
				4'b0001:out[7:0]=8'b10011111;
				4'b0010:out[7:0]=8'b00100101;
				4'b0011:out[7:0]=8'b00001101;
				4'b0100:out[7:0]=8'b10011001;
				4'b0101:out[7:0]=8'b01001001;
				4'b0110:out[7:0]=8'b01000001;
				4'b0111:out[7:0]=8'b00011111;
				4'b1000:out[7:0]=8'b00000001;
				4'b1001:out[7:0]=8'b00001001;
				4'b1010:out[7:0]=8'b00010001;
				4'b1011:out[7:0]=8'b11000001;
				4'b1100:out[7:0]=8'b01100011;
				4'b1101:out[7:0]=8'b10000101;
				4'b1110:out[7:0]=8'b01100001;
				4'b1111:out[7:0]=8'b01110001;
			endcase

			case(in[7:4])
				4'b0000:out[15:8]=8'b00000011;
				4'b0001:out[15:8]=8'b10011111;
				4'b0010:out[15:8]=8'b00100101;
				4'b0011:out[15:8]=8'b00001101;
				4'b0100:out[15:8]=8'b10011001;
				4'b0101:out[15:8]=8'b01001001;
				4'b0110:out[15:8]=8'b01000001;
				4'b0111:out[15:8]=8'b00011111;
				4'b1000:out[15:8]=8'b00000001;
				4'b1001:out[15:8]=8'b00001001;
				4'b1010:out[15:8]=8'b00010001;
				4'b1011:out[15:8]=8'b11000001;
				4'b1100:out[15:8]=8'b01100011;
				4'b1101:out[15:8]=8'b10000101;
				4'b1110:out[15:8]=8'b01100001;
				4'b1111:out[15:8]=8'b01110001;
			endcase

			case(in[11:8])
				4'b0000:out[23:16]=8'b00000011;
				4'b0001:out[23:16]=8'b10011111;
				4'b0010:out[23:16]=8'b00100101;
				4'b0011:out[23:16]=8'b00001101;
				4'b0100:out[23:16]=8'b10011001;
				4'b0101:out[23:16]=8'b01001001;
				4'b0110:out[23:16]=8'b01000001;
				4'b0111:out[23:16]=8'b00011111;
				4'b1000:out[23:16]=8'b00000001;
				4'b1001:out[23:16]=8'b00001001;
				4'b1010:out[23:16]=8'b00010001;
				4'b1011:out[23:16]=8'b11000001;
				4'b1100:out[23:16]=8'b01100011;
				4'b1101:out[23:16]=8'b10000101;
				4'b1110:out[23:16]=8'b01100001;
				4'b1111:out[23:16]=8'b01110001;
			endcase

			case(in[15:12])
				4'b0000:out[31:24]=8'b00000011;
				4'b0001:out[31:24]=8'b10011111;
				4'b0010:out[31:24]=8'b00100101;
				4'b0011:out[31:24]=8'b00001101;
				4'b0100:out[31:24]=8'b10011001;
				4'b0101:out[31:24]=8'b01001001;
				4'b0110:out[31:24]=8'b01000001;
				4'b0111:out[31:24]=8'b00011111;
				4'b1000:out[31:24]=8'b00000001;
				4'b1001:out[31:24]=8'b00001001;
				4'b1010:out[31:24]=8'b00010001;
				4'b1011:out[31:24]=8'b11000001;
				4'b1100:out[31:24]=8'b01100011;
				4'b1101:out[31:24]=8'b10000101;
				4'b1110:out[31:24]=8'b01100001;
				4'b1111:out[31:24]=8'b01110001;
			endcase

			case(in[19:16])
				4'b0000:out[39:32]=8'b00000011;
				4'b0001:out[39:32]=8'b10011111;
				4'b0010:out[39:32]=8'b00100101;
				4'b0011:out[39:32]=8'b00001101;
				4'b0100:out[39:32]=8'b10011001;
				4'b0101:out[39:32]=8'b01001001;
				4'b0110:out[39:32]=8'b01000001;
				4'b0111:out[39:32]=8'b00011111;
				4'b1000:out[39:32]=8'b00000001;
				4'b1001:out[39:32]=8'b00001001;
				4'b1010:out[39:32]=8'b00010001;
				4'b1011:out[39:32]=8'b11000001;
				4'b1100:out[39:32]=8'b01100011;
				4'b1101:out[39:32]=8'b10000101;
				4'b1110:out[39:32]=8'b01100001;
				4'b1111:out[39:32]=8'b01110001;
			endcase

			case(in[23:20])
				4'b0000:out[47:40]=8'b00000011;
				4'b0001:out[47:40]=8'b10011111;
				4'b0010:out[47:40]=8'b00100101;
				4'b0011:out[47:40]=8'b00001101;
				4'b0100:out[47:40]=8'b10011001;
				4'b0101:out[47:40]=8'b01001001;
				4'b0110:out[47:40]=8'b01000001;
				4'b0111:out[47:40]=8'b00011111;
				4'b1000:out[47:40]=8'b00000001;
				4'b1001:out[47:40]=8'b00001001;
				4'b1010:out[47:40]=8'b00010001;
				4'b1011:out[47:40]=8'b11000001;
				4'b1100:out[47:40]=8'b01100011;
				4'b1101:out[47:40]=8'b10000101;
				4'b1110:out[47:40]=8'b01100001;
				4'b1111:out[47:40]=8'b01110001;
			endcase

			case(in[27:24])
				4'b0000:out[55:48]=8'b00000011;
				4'b0001:out[55:48]=8'b10011111;
				4'b0010:out[55:48]=8'b00100101;
				4'b0011:out[55:48]=8'b00001101;
				4'b0100:out[55:48]=8'b10011001;
				4'b0101:out[55:48]=8'b01001001;
				4'b0110:out[55:48]=8'b01000001;
				4'b0111:out[55:48]=8'b00011111;
				4'b1000:out[55:48]=8'b00000001;
				4'b1001:out[55:48]=8'b00001001;
				4'b1010:out[55:48]=8'b00010001;
				4'b1011:out[55:48]=8'b11000001;
				4'b1100:out[55:48]=8'b01100011;
				4'b1101:out[55:48]=8'b10000101;
				4'b1110:out[55:48]=8'b01100001;
				4'b1111:out[55:48]=8'b01110001;
			endcase

			case(in[31:28])
				4'b0000:out[63:56]=8'b00000011;
				4'b0001:out[63:56]=8'b10011111;
				4'b0010:out[63:56]=8'b00100101;
				4'b0011:out[63:56]=8'b00001101;
				4'b0100:out[63:56]=8'b10011001;
				4'b0101:out[63:56]=8'b01001001;
				4'b0110:out[63:56]=8'b01000001;
				4'b0111:out[63:56]=8'b00011111;
				4'b1000:out[63:56]=8'b00000001;
				4'b1001:out[63:56]=8'b00001001;
				4'b1010:out[63:56]=8'b00010001;
				4'b1011:out[63:56]=8'b11000001;
				4'b1100:out[63:56]=8'b01100011;
				4'b1101:out[63:56]=8'b10000101;
				4'b1110:out[63:56]=8'b01100001;
				4'b1111:out[63:56]=8'b01110001;
			endcase


	end
endmodule
